interface shift_reg_intf;
    bit       d;
    bit       clk;
    bit       en;
    bit       dir;
    bit       rstn;
    bit [7:0] out;
endinterface : shift_reg_intf
